module fadd32_tb;
endmodule