// Author: Ninaad Desai
// Description: 24-bit barrel logical right shifter with even rounding-off  
module sr24(
    input [23:0] oprnd,
    input [4:0] shamt,
    output [23:0] reslt
);
endmodule