module comp8_tb;
    reg [7:0] a;
    reg [7:0] b;
endmodule